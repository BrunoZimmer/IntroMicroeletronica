* SPICE NETLIST
***************************************

.SUBCKT CELL A B C Gnd Vdd Y
** N=9 EP=6 IP=0 FDC=8
M0 4 A 5 Gnd NMOS_VTL L=5e-08 W=3e-07 AD=6.45e-14 AS=8.55e-14 PD=1.03e-06 PS=1.17e-06 $X=164895 $Y=81225 $D=1
M1 5 B 4 Gnd NMOS_VTL L=5e-08 W=3e-07 AD=1.155e-13 AS=6.45e-14 PD=1.37e-06 PS=1.03e-06 $X=165425 $Y=81225 $D=1
M2 Gnd C 5 Gnd NMOS_VTL L=5e-08 W=3e-07 AD=6.975e-14 AS=1.155e-13 PD=1.065e-06 PS=1.37e-06 $X=166295 $Y=81225 $D=1
M3 Y 4 Gnd Gnd NMOS_VTL L=5e-08 W=3e-07 AD=5.7e-14 AS=6.975e-14 PD=9.8e-07 PS=1.065e-06 $X=166860 $Y=81225 $D=1
M4 2 A Vdd Vdd PMOS_VTL L=5e-08 W=6e-07 AD=1.29e-13 AS=1.71e-13 PD=1.63e-06 PS=1.77e-06 $X=164895 $Y=83465 $D=0
M5 4 B 2 Vdd PMOS_VTL L=5e-08 W=6e-07 AD=2.31e-13 AS=1.29e-13 PD=1.97e-06 PS=1.63e-06 $X=165425 $Y=83465 $D=0
M6 Vdd C 4 Vdd PMOS_VTL L=5e-08 W=6e-07 AD=1.395e-13 AS=2.31e-13 PD=1.665e-06 PS=1.97e-06 $X=166295 $Y=83465 $D=0
M7 Y 4 Vdd Vdd PMOS_VTL L=5e-08 W=6e-07 AD=1.05e-13 AS=1.395e-13 PD=1.55e-06 PS=1.665e-06 $X=166860 $Y=83465 $D=0
.ENDS
***************************************

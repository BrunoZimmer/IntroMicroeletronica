*Tristate non-inverter

.SUBCKT TNI IN ZN EN ENB VDD VSS 
*M_i Drain Gate Source Bulk
M_i_0 1 IN VSS VSS NMOS W=0.415000U L=0.050000U
M_i_2 ZN ENB 1 VSS NMOS W=0.415000U L=0.050000U

M_i_3 ZN EN 2 VDD PMOS W=0.630000U L=0.050000U
M_i_1 2 IN VDD VDD PMOS W=0.630000U L=0.050000U

.ENDS 

